 -- 
 -- Copyright (c) 2023, Daniel Lammers, Amir Moradi, Nicolai Müller, Aein Rezaei Shahmirzadi
 -- 
 -- All rights reserved.
 -- 
 -- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
 -- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
 -- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
 -- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
 -- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
 -- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
 -- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
 -- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
 -- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
 -- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
 -- 
 -- Please see LICENSE and README for license and further instructions.
 -- 

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

entity TB_RAMBAM_AES is
end TB_RAMBAM_AES;

architecture Behavioral of TB_RAMBAM_AES is

	component Circuit is
		Generic ( d    : integer := 8;
					 n    : integer := 8;
					 m    : integer := 8;
					 Mul2 : std_logic_vector := "0001011000000000100010110000000001000101000000000011010000000000000110100000000010011011000000000101101100000000001011010000000000000000000101100000000010001011000000000100010100000000001101000000000000011010000000001001101100000000010110110000000000101101";
				    Mul3 : std_logic_vector := "1001011000000000110010110000000001100101000000000010010000000000000100100000000010011111000000000101100100000000001011000000000000000000100101100000000011001011000000000110010100000000001001000000000000010010000000001001111100000000010110010000000000101100";
					 RInv : std_logic_vector := "1011001101101011001110000010101101110110000000110001100100010001";
					 R    : std_logic_vector := "1010011101010000000101110011010000000011010010100011000100110101";
					 TInv : std_logic_vector := "1001010011001010111001010110011000110011100011010101001000101001";
					 T    : std_logic_vector := "1011110101011110001011111010101001010101100101111111011001111011";
					 poly : std_logic_vector := "10000000000000011";
					 A    : std_logic_vector := "0000001000000000000010010000000011111110000000000011111100000000001010010000000000010001000000000110010000000000011010010000000000000000111011010000000000111111000000000000010000000000010010110000000000100001000000000111100100000000000000100000000000001100";
					 Q0	: std_logic_vector := "1000111000000000000000110000000001000111000000000000111100000000001000000000000000001001000000000001110100000000000001110000000000000000111010000000000000111000000000000111010000000000111101000000000000000010000000001001001000000000110100010000000001110001";
					 Q1	: std_logic_vector := "1011101000000000000110100000000000010000000000000011001100000000010001110000000000100111000000000010000100000000000100110000000000000000101001100000000010000010000000000010101000000000110000100000000011010001000000001100110100000000010101010000000011001001";
					 Q3	: std_logic_vector := "1111111100000000010101010000000000110011000000000001000100000000000011110000000000000101000000000000001100000000000000010000000000000000000101000000000011110011000000001010111000000000011100010000000000101111000000001111000100000000010001000000000000111100";
					 C	   : std_logic_vector := x"009b");
		Port ( clk 	      : in  std_logic;
				 rst 	      : in  std_logic;
				 en			: in  std_logic;
				 en_in      : in  std_logic;
				 en_out     : in  std_logic;
				 x0 		   : in  std_logic_vector(127 downto 0);
			    x1 		   : in  std_logic_vector(127 downto 0);
				 key0 	   : in  std_logic_vector(127 downto 0);
			    key1 	   : in  std_logic_vector(127 downto 0);
				
				 randomness : in  std_logic_vector(1119 downto 0); -- 8*7*(16+4)
				
				 done       : out std_logic;
			    z0 		   : out std_logic_vector(127 downto 0);
			    z1 		   : out std_logic_vector(127 downto 0));
	end component;

	signal   clk        : std_logic;
	constant clk_period : time := 10 ns;
	
	signal x0, x1, key0, key1, z0, z1 : std_logic_vector(127 downto 0);

	signal randomness_reshares : std_logic_vector(1119 downto 0);
	
	signal en, en_in, en_out, rst, done : std_logic;

begin

   uut: Circuit
		generic map (
			d    => 8,
			n    => 8,
			m    => 8,
			Mul2 => "0001011000000000100010110000000001000101000000000011010000000000000110100000000010011011000000000101101100000000001011010000000000000000000101100000000010001011000000000100010100000000001101000000000000011010000000001001101100000000010110110000000000101101",
			Mul3 => "1001011000000000110010110000000001100101000000000010010000000000000100100000000010011111000000000101100100000000001011000000000000000000100101100000000011001011000000000110010100000000001001000000000000010010000000001001111100000000010110010000000000101100",
			RInv => "1011001101101011001110000010101101110110000000110001100100010001",
			R    => "1010011101010000000101110011010000000011010010100011000100110101",
			TInv => "1001010011001010111001010110011000110011100011010101001000101001",
			T    => "1011110101011110001011111010101001010101100101111111011001111011",
			poly => "10000000000000011",
			A    => "0000001000000000000010010000000011111110000000000011111100000000001010010000000000010001000000000110010000000000011010010000000000000000111011010000000000111111000000000000010000000000010010110000000000100001000000000111100100000000000000100000000000001100",
		   Q0	  => "1000111000000000000000110000000001000111000000000000111100000000001000000000000000001001000000000001110100000000000001110000000000000000111010000000000000111000000000000111010000000000111101000000000000000010000000001001001000000000110100010000000001110001",
		   Q1	  => "1011101000000000000110100000000000010000000000000011001100000000010001110000000000100111000000000010000100000000000100110000000000000000101001100000000010000010000000000010101000000000110000100000000011010001000000001100110100000000010101010000000011001001",
		   Q3	  => "1111111100000000010101010000000000110011000000000001000100000000000011110000000000000101000000000000001100000000000000010000000000000000000101000000000011110011000000001010111000000000011100010000000000101111000000001111000100000000010001000000000000111100",
		   C	  => x"009b"
		)
		port map (
			clk 	     => clk,
			rst 	     => rst,
			en			  => en,
			en_in      => en_in,
			en_out     => en_out,
			x0 	     => x0,
			x1 	     => x1,
			key0       => key0,
			key1       => key1,

		   randomness => randomness_reshares,

			done       => done,
			z0 	     => z0,
			z1 	     => z1
		);		
		
	clk_process: process
	begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
	end process;

	stim_proc: process
   begin			
		en  <= '0';
		rst <= '1';
		
		wait for clk_period;
		
		-- inputs can change here --
		x0 <= x"0895db6dba58e0df9e9a88acd4d2405b";
		x1 <= x"00000000000000000000000000000000";
		
		key0 <= x"e696f30db27608f20a07f92a1c37fff4";
		key1 <= x"00000000000000000000000000000000";
		
		randomness_reshares <= x"e60b675d938dfbef323bd4e58ef0aacabc6787881030b80668ea72943ac9008d005e03c18e0003ead7ab974a9a371ef28b17036f7689ed1345a79e60b75e2e3a423926d4a48e02445341fd4baa38e4d6621b5997c550fc9ab59f3b8f1a79e0c6ec9839472a4a786a9c1167c1d8f9d9845a46cf7cc311114b3182c60360a72aafc7e9e57b01d52d55766dd691";--(others => '0');
		-- ---------------------- --
		
		rst <= '0';
		
		wait for clk_period;
		
		en_in <= '1';
		
		wait for clk_period;
		
		en_in <= '0';      
		en  <= '1';
		
		wait until (done = '1');
		
		wait for clk_period;
		
		en_out <= '1';
		
		wait for clk_period;
		
		en_out <= '0';
		
		assert((z0 xor z1) = x"0573702ebc4fdabd750830903cc554c6")
	    report "error" severity failure; 

      wait;
   end process;

end Behavioral;

